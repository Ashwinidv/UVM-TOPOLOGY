/////-----------------------------------------------------------------------------------------------////
////----------------------------------UVM_PACKAGE---------------------------------------------------////
////------------------------------------------------------------------------------------------------////

   
  
package basic_pkg;
   import uvm_pkg::*;

   
  `include "uvm_sequence_item.sv"
  `include "uvm_sequence.sv"
  `include "uvm_sequencer.sv"
  `include "uvm_driver.sv"
  `include "uvm_monitor.sv"
  `include "uvm_agent.sv"
  `include "uvm_scoreboard.sv"
  `include "uvm_env.sv"
  `include "uvm_test.sv"


endpackage : basic_pkg
